module BRAMDSP(
    CLK1, CLK2,
    A1ADDR, A2ADDR, A1EN, A2EN, A1DATA, A2DATA,
    B1ADDR, B2ADDR, B3ADDR, B4ADDR, B1EN, B2EN, B3EN, B4EN, B1DATA, B2DATA, B3DATA, B4DATA,
    C1ADDR, C2ADDR, C3ADDR, C4ADDR, C1EN, C2EN, C3EN, C4EN, C1DATA, C2DATA, C3DATA, C4DATA);

parameter CFG_ABITS = 11;
parameter CFG_DBITS = 32;
parameter CFG_ENABLE_A = 2;
parameter CFG_ENABLE_B = 4;
parameter CFG_ENABLE_C = 4;

input CLK1, CLK2;
input [CFG_ABITS-1:0] A1ADDR, A2ADDR, B1ADDR, B2ADDR, B3ADDR, B4ADDR, C1ADDR, C2ADDR, C3ADDR, C4ADDR;
output [CFG_DBITS-1:0] A1DATA, A2DATA;
input [CFG_DBITS-1:0] B1DATA, B2DATA, B3DATA, B4DATA;
input [CFG_DBITS-1:0] C1DATA, C2DATA, C3DATA, C4DATA;
input [CFG_ENABLE_A-1:0] A1EN, A2EN;
input [CFG_ENABLE_B-1:0] B1EN, B2EN, B3EN, B4EN;
input [CFG_ENABLE_C-1:0] C1EN, C2EN, C3EN, C4EN;

endmodule